// Benchmark "c432_default" written by ABC on Mon Dec 01 21:12:31 2025

module c432_default ( 
    in4, in17, in30, in43, in56, in69, in82, in95, in108, in1, in11, in24,
    in37, in50, in63, in76, in89, in102, in8, in21, in34, in47, in60, in73,
    in86, in99, in112, in14, in27, in40, in53, in66, in79, in92, in105,
    in115,
    out223, out329, out370, out421, out430, out431, out432  );
  input  in4, in17, in30, in43, in56, in69, in82, in95, in108, in1, in11,
    in24, in37, in50, in63, in76, in89, in102, in8, in21, in34, in47, in60,
    in73, in86, in99, in112, in14, in27, in40, in53, in66, in79, in92,
    in105, in115;
  output out223, out329, out370, out421, out430, out431, out432;
  wire n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n98, n99,
    n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n293, n294,
    n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
    n308, n309, n310, n311, n312, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323;
  assign n43 = ~in108;
  assign n44 = ~in1;
  assign n45 = ~in11;
  assign n46 = ~in24;
  assign n47 = ~in37;
  assign n48 = ~in50;
  assign n49 = ~in63;
  assign n50 = ~in76;
  assign n51 = ~in89;
  assign n52 = ~in102;
  assign n53 = ~in8;
  assign n54 = ~in21;
  assign n55 = ~in34;
  assign n56 = ~in47;
  assign n57 = ~in60;
  assign n58 = ~in73;
  assign n59 = ~in86;
  assign n60 = ~in99;
  assign n61 = ~in112;
  assign n62 = ~in14;
  assign n63 = ~in27;
  assign n64 = ~in40;
  assign n65 = ~in53;
  assign n66 = ~in66;
  assign n67 = ~in79;
  assign n68 = ~in92;
  assign n69 = ~in105;
  assign n70 = ~in115;
  assign n71 = in56 & n48;
  assign n72 = ~n71;
  assign n73 = in30 & n46;
  assign n74 = ~n73;
  assign n75 = in17 & n45;
  assign n76 = ~n75;
  assign n77 = n74 & n76;
  assign n78 = in69 & n49;
  assign n79 = ~n78;
  assign n80 = in43 & n47;
  assign n81 = ~n80;
  assign n82 = n79 & n81;
  assign n83 = n77 & n82;
  assign n84 = n72 & n83;
  assign n85 = in108 & n52;
  assign n86 = ~n85;
  assign n87 = in4 & n44;
  assign n88 = ~n87;
  assign n89 = n86 & n88;
  assign n90 = in95 & n51;
  assign n91 = ~n90;
  assign n92 = in82 & n50;
  assign n93 = ~n92;
  assign n94 = n91 & n93;
  assign n95 = n89 & n94;
  assign n96 = n84 & n95;
  assign out223 = ~n96;
  assign n98 = n81 & out223;
  assign n99 = ~n98;
  assign n100 = n56 & n99;
  assign n101 = in43 & n100;
  assign n102 = ~n101;
  assign n103 = n72 & out223;
  assign n104 = ~n103;
  assign n105 = n57 & n104;
  assign n106 = in56 & n105;
  assign n107 = ~n106;
  assign n108 = n102 & n107;
  assign n109 = n79 & out223;
  assign n110 = ~n109;
  assign n111 = n58 & n110;
  assign n112 = in69 & n111;
  assign n113 = ~n112;
  assign n114 = n93 & out223;
  assign n115 = ~n114;
  assign n116 = n59 & n115;
  assign n117 = in82 & n116;
  assign n118 = ~n117;
  assign n119 = n113 & n118;
  assign n120 = n88 & out223;
  assign n121 = ~n120;
  assign n122 = n53 & n121;
  assign n123 = in4 & n122;
  assign n124 = ~n123;
  assign n125 = n74 & out223;
  assign n126 = ~n125;
  assign n127 = n55 & n126;
  assign n128 = ~n127;
  assign n129 = in30 & n127;
  assign n130 = ~n129;
  assign n131 = n76 & out223;
  assign n132 = ~n131;
  assign n133 = n54 & n132;
  assign n134 = ~n133;
  assign n135 = in17 & n133;
  assign n136 = ~n135;
  assign n137 = n130 & n136;
  assign n138 = n124 & n137;
  assign n139 = n91 & out223;
  assign n140 = ~n139;
  assign n141 = n60 & n140;
  assign n142 = in95 & n141;
  assign n143 = ~n142;
  assign n144 = n86 & out223;
  assign n145 = ~n144;
  assign n146 = n61 & n145;
  assign n147 = in108 & n146;
  assign n148 = ~n147;
  assign n149 = n143 & n148;
  assign n150 = n138 & n149;
  assign n151 = n119 & n150;
  assign n152 = n108 & n151;
  assign out329 = ~n152;
  assign n154 = n66 & n104;
  assign n155 = n107 & out329;
  assign n156 = ~n155;
  assign n157 = in56 & n156;
  assign n158 = n154 & n157;
  assign n159 = ~n158;
  assign n160 = n134 & out329;
  assign n161 = ~n160;
  assign n162 = in17 & n161;
  assign n163 = n63 & n132;
  assign n164 = n162 & n163;
  assign n165 = ~n164;
  assign n166 = n64 & n126;
  assign n167 = n128 & out329;
  assign n168 = ~n167;
  assign n169 = in30 & n168;
  assign n170 = n166 & n169;
  assign n171 = ~n170;
  assign n172 = n165 & n171;
  assign n173 = n67 & n110;
  assign n174 = n113 & out329;
  assign n175 = ~n174;
  assign n176 = in69 & n175;
  assign n177 = n173 & n176;
  assign n178 = ~n177;
  assign n179 = n102 & out329;
  assign n180 = ~n179;
  assign n181 = n65 & n99;
  assign n182 = in43 & n181;
  assign n183 = n180 & n182;
  assign n184 = ~n183;
  assign n185 = n178 & n184;
  assign n186 = n172 & n185;
  assign n187 = n159 & n186;
  assign n188 = n62 & n121;
  assign n189 = n124 & out329;
  assign n190 = ~n189;
  assign n191 = in4 & n190;
  assign n192 = n188 & n191;
  assign n193 = ~n192;
  assign n194 = n148 & out329;
  assign n195 = ~n194;
  assign n196 = in108 & n195;
  assign n197 = n70 & n145;
  assign n198 = n196 & n197;
  assign n199 = ~n198;
  assign n200 = n193 & n199;
  assign n201 = n69 & n140;
  assign n202 = n143 & out329;
  assign n203 = ~n202;
  assign n204 = in95 & n203;
  assign n205 = n201 & n204;
  assign n206 = ~n205;
  assign n207 = n118 & out329;
  assign n208 = ~n207;
  assign n209 = in82 & n208;
  assign n210 = n68 & n115;
  assign n211 = n209 & n210;
  assign n212 = ~n211;
  assign n213 = n206 & n212;
  assign n214 = n200 & n213;
  assign n215 = n187 & n214;
  assign out370 = ~n215;
  assign n217 = in99 & out329;
  assign n218 = ~n217;
  assign n219 = in105 & out370;
  assign n220 = ~n219;
  assign n221 = n218 & n220;
  assign n222 = in89 & out223;
  assign n223 = ~n222;
  assign n224 = in95 & n223;
  assign n225 = n221 & n224;
  assign n226 = ~n225;
  assign n227 = in92 & out370;
  assign n228 = ~n227;
  assign n229 = in86 & out329;
  assign n230 = ~n229;
  assign n231 = n228 & n230;
  assign n232 = in76 & out223;
  assign n233 = ~n232;
  assign n234 = in82 & n233;
  assign n235 = n231 & n234;
  assign n236 = ~n235;
  assign n237 = in63 & out223;
  assign n238 = ~n237;
  assign n239 = in69 & n238;
  assign n240 = in79 & out370;
  assign n241 = ~n240;
  assign n242 = in73 & out329;
  assign n243 = ~n242;
  assign n244 = n241 & n243;
  assign n245 = n239 & n244;
  assign n246 = ~n245;
  assign n247 = n236 & n246;
  assign n248 = ~n247;
  assign n249 = in37 & out223;
  assign n250 = ~n249;
  assign n251 = in43 & n250;
  assign n252 = in47 & out329;
  assign n253 = ~n252;
  assign n254 = in53 & out370;
  assign n255 = ~n254;
  assign n256 = n253 & n255;
  assign n257 = n251 & n256;
  assign n258 = ~n257;
  assign n259 = in24 & out223;
  assign n260 = ~n259;
  assign n261 = in30 & n260;
  assign n262 = in34 & out329;
  assign n263 = ~n262;
  assign n264 = in40 & out370;
  assign n265 = ~n264;
  assign n266 = n263 & n265;
  assign n267 = n261 & n266;
  assign n268 = ~n267;
  assign n269 = in11 & out223;
  assign n270 = ~n269;
  assign n271 = in17 & n270;
  assign n272 = in21 & out329;
  assign n273 = ~n272;
  assign n274 = in27 & out370;
  assign n275 = ~n274;
  assign n276 = n273 & n275;
  assign n277 = n271 & n276;
  assign n278 = ~n277;
  assign n279 = in50 & out223;
  assign n280 = ~n279;
  assign n281 = in56 & n280;
  assign n282 = in60 & out329;
  assign n283 = ~n282;
  assign n284 = in66 & out370;
  assign n285 = ~n284;
  assign n286 = n283 & n285;
  assign n287 = n281 & n286;
  assign n288 = ~n287;
  assign n289 = n278 & n288;
  assign n290 = n268 & n289;
  assign n291 = n258 & n290;
  assign out430 = ~n291;
  assign n293 = n247 & n291;
  assign n294 = n43 & n293;
  assign n295 = n226 & n294;
  assign n296 = ~n295;
  assign n297 = in8 & out329;
  assign n298 = ~n297;
  assign n299 = in4 & n298;
  assign n300 = in14 & out370;
  assign n301 = ~n300;
  assign n302 = in1 & out223;
  assign n303 = ~n302;
  assign n304 = n301 & n303;
  assign n305 = n299 & n304;
  assign n306 = ~n305;
  assign out421 = n296 & n306;
  assign n308 = n248 & n258;
  assign n309 = n288 & n308;
  assign n310 = ~n309;
  assign n311 = n278 & n310;
  assign n312 = n268 & n311;
  assign out431 = ~n312;
  assign n314 = n236 & n225;
  assign n315 = ~n314;
  assign n316 = n245 & n288;
  assign n317 = ~n316;
  assign n318 = n315 & n317;
  assign n319 = n258 & n318;
  assign n320 = ~n319;
  assign n321 = n268 & n320;
  assign n322 = ~n321;
  assign n323 = n278 & n322;
  assign out432 = ~n323;
endmodule


